** Profile: "BitTest-stdBitSliceTest"  [ C:\Users\Joe2TB\Documents\ECE424\OrCAD\PCB_Assign2-PSpiceFiles\BitTest\stdBitSliceTest.sim ] 

** Creating circuit file "stdBitSliceTest.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.STMLIB "../../../pcb_assign2-pspicefiles/pcb_assign2.stl" 
* From [PSPICE NETLIST] section of C:\Users\Joe2TB\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\BitTest.net" 


.END
